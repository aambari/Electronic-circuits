Fatal Error: Previous analysis already found: .tran 50us 2ms
