BASIC_AMPLIFIER.CIR - DISCRETE AMPLIFIER
*
VS	1	0	AC 1	SIN(0 0.1V 1KHZ)
CIN	1	2	1UF
RIN1	2	0	100K
*
* POWER SUPPLIES
VCC	100	0	DC	+15V
VEE	101	0	DC	-15V
* 
* DIFF AMP
RE	100	8	14.3K
Q1	4 2 	8	QPNP
Q2	101 3	8	QPNP
RC1	4	101	1800
*
* GAIN STAGE AND COMPENSATION
Q3	14 4	101	QNPN3
CC	14	4	10PF
*
* OUTPUT STAGE BIAS
RC3	100	11	4K
D1	11	13	D1N4148
D2	13	14	D1N4148
*
* OUTPUT STAGE
Q4	100 11	20	QNPN4
Q5	101 14	20	QPNP5
*
* LOAD
RL	20	0	100000
*
* FEEDBACK
RF2	20	3	100K
RF1	3	21	11K
CF1	21	0	10UF
*
* SMALL SIGNAL DEVICES
.model	QNPN	NPN(BF=100)
.model	QPNP	PNP(BF=100)
.model	QNPN3	NPN(BF=100)
.model	D1N4148	D(Is=0.1p Rs=16 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

* OUTPUT POWER DEVICES
.model	QNPN4	NPN(BF=100)
.model	QPNP5	PNP(BF=100)

*
.TRAN	50US 2MS
.AC DEC 5 1 1MEG
.PROBE
.END